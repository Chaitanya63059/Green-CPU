`timescale 1ns / 1ps

module mux2 #(parameter WIDTH = 16)(
    input  [WIDTH-1:0] d0, d1,
    input               sel,
    output [WIDTH-1:0] y
);



endmodule