`timescale 1ns / 1ps

module mux3 #(parameter WIDTH = 16)(
    input       [15:0] d0, d1, d2,
    input       [1:0] sel,
    output      [15:0] y
);


endmodule

