`timescale 1ns / 1ps

// adder.v - logic for adder

module adder #(parameter WIDTH = 16) (
    input       [WIDTH-1:0] a, b,
    output      [WIDTH-1:0] sum
);



endmodule

